class ahbl_mst_sqr extends uvm_sequencer #(ahbl_tran);
  `uvm_component_utils(ahbl_mst_sqr)

  function new(string name, uvm_component parent);
    super.new(name,parent);
  endfunction

endclass
