`ifndef TEST_LIB_SV
`define TEST_LIB_SV

`include "./ahbl_mst_single_read32.sv"
`include "./ahbl_mst_single_write32_apb_slv_nrdy.sv"
`include "./ahbl_mst_burst.sv"
`include "./ahbl_mst_burst_apb_slv_slverr.sv"
`include "./ahbl_mst_tight_transfer.sv"

`endif
