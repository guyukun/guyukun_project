package ahb2apb_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  
  import apb_slv_pkg::*;
  import ahbl_mst_pkg::*;

  `include "func_cov.sv"
  `include "ahb2apb_scb.sv"
  `include "ahb2apb_env.sv"
endpackage
